module bindfiles;
	bind ammon_lc3 lc3_asserts p1 (.*);
endmodule
